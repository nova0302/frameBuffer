//                            -*- Mode: Verilog -*-
//
// Filename: defines.sv
// Created: Sun Feb  8 12:28:49 2015 (+0900)
// Last-Updated:
//           By:
//     Update #: 3

//
// defines.sv ends here
`define SIMULATION
